module mux6_test();
	



endmodule 