module deco1(input logic[2:0] color_in, 
			output logic [23:0]color_out);

	logic[23:0] color_out_temp;
	
	assign color_out = {color_out_temp[7:0], color_out_temp[15:8], color_out_temp[23:16]};
	
	always_comb
		case(color_in)
			3'd0:color_out_temp = 24'h000000;
			3'd1:color_out_temp = 24'h000000;
			3'd2:color_out_temp = 24'h00fff0;
			3'd3:color_out_temp = 24'hffffff;
			3'd4:color_out_temp = 24'h0087ff;
			default : color_out_temp = 24'h0;
		endcase


/* Piskel data for "Flappy" */
/* 0x00000000=0   
 * 0xff000000=1
 * 0xff00fff0=2
 * 0xffffffff=3
 * 4=0xff0087ff
 * */
		
endmodule 