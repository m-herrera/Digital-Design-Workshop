module overflow_flag_test();



endmodule 